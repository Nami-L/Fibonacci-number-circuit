`timescale 1ns/1ps

package fsm_fino_pkg;
// Define the state for the Fibonacci number fsm_fino_pkg

typedef enum {
    IDLE,
    OP,
    DONE,
    XXX // Uundefined states
}state_e;

endpackage: fsm_fino_pkg



